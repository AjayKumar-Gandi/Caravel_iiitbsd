* NGSPICE file created from iiitb_sdm.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

.subckt iiitb_sdm clock detector_out reset sequence_in vccd1 vssd1
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_29_ input1/X _29_/D vssd1 vssd1 vccd1 vccd1 _29_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__23__A _28_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_28_ _28_/A vssd1 vssd1 vccd1 vccd1 _28_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27_ _28_/A vssd1 vssd1 vccd1 vccd1 _27_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26_ _26_/A vssd1 vssd1 vccd1 vccd1 _29_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25_ _32_/Q _25_/B _25_/C vssd1 vssd1 vccd1 vccd1 _26_/A sky130_fd_sc_hd__and3_1
XFILLER_38_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24_ _31_/Q _30_/Q _24_/C vssd1 vssd1 vccd1 vccd1 _25_/C sky130_fd_sc_hd__and3b_1
XFILLER_37_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__29__D _29_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23_ _28_/A vssd1 vssd1 vccd1 vccd1 _25_/B sky130_fd_sc_hd__inv_2
XFILLER_187_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22_ _20_/Y _30_/Q _14_/B _18_/B _21_/X vssd1 vssd1 vccd1 vccd1 _32_/D sky130_fd_sc_hd__o2111a_1
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__31__CLK input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_6587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21_ _31_/Q _32_/Q vssd1 vssd1 vccd1 vccd1 _21_/X sky130_fd_sc_hd__or2_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20_ _31_/Q vssd1 vssd1 vccd1 vccd1 _20_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput1 clock vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_8
XFILLER_211_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1022 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput2 reset vssd1 vssd1 vccd1 vccd1 _28_/A sky130_fd_sc_hd__buf_4
XFILLER_83_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1034 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput3 sequence_in vssd1 vssd1 vccd1 vccd1 _24_/C sky130_fd_sc_hd__buf_6
XFILLER_84_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1046 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16__B _24_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__27__A _28_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_7059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__24__C _24_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__30__CLK input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19_ _19_/A vssd1 vssd1 vccd1 vccd1 _31_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18_ _32_/Q _18_/B _18_/C vssd1 vssd1 vccd1 vccd1 _19_/A sky130_fd_sc_hd__and3b_1
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17_ _31_/Q _30_/Q vssd1 vssd1 vccd1 vccd1 _18_/C sky130_fd_sc_hd__xor2_1
XFILLER_93_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1031 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16_ _30_/Q _24_/C vssd1 vssd1 vccd1 vccd1 _18_/B sky130_fd_sc_hd__xor2_1
XFILLER_53_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_32_ input1/X _32_/D _28_/Y vssd1 vssd1 vccd1 vccd1 _32_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15_ _15_/A vssd1 vssd1 vccd1 vccd1 _30_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_7152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1003 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14__A _24_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_31_ input1/X _31_/D _27_/Y vssd1 vssd1 vccd1 vccd1 _31_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14_ _24_/C _14_/B vssd1 vssd1 vccd1 vccd1 _15_/A sky130_fd_sc_hd__and2_1
XFILLER_4_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_30_ input1/X _30_/D _25_/B vssd1 vssd1 vccd1 vccd1 _30_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13_ _31_/Q _32_/Q vssd1 vssd1 vccd1 vccd1 _14_/B sky130_fd_sc_hd__nand2_1
XFILLER_187_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__28__A _28_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_A sequence_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__29__CLK input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input1_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput4 _29_/Q vssd1 vssd1 vccd1 vccd1 detector_out sky130_fd_sc_hd__buf_2
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_7138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1721 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_7661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1777 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_7491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_1353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1917 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__32__CLK input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1665 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1789 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
.ends

