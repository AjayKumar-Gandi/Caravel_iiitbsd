magic
tech sky130B
magscale 1 2
timestamp 1662965546
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 14 2128 179754 117552
<< metal2 >>
rect 32862 119200 32918 120000
rect 179694 119200 179750 120000
rect 18 0 74 800
rect 146850 0 146906 800
<< obsm2 >>
rect 20 119144 32806 119354
rect 32974 119144 179638 119354
rect 20 856 179748 119144
rect 130 800 146794 856
rect 146962 800 179748 856
<< obsm3 >>
rect 4210 2143 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 18 0 74 800 6 clock
port 1 nsew signal input
rlabel metal2 s 32862 119200 32918 120000 6 detector_out
port 2 nsew signal output
rlabel metal2 s 179694 119200 179750 120000 6 reset
port 3 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 sequence_in
port 4 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5503798
string GDS_FILE /home/ajaykumar/Desktop/Caravel_iiitbsd/openlane/iiitb_sdm/runs/22_09_12_12_17/results/signoff/iiitb_sdm.magic.gds
string GDS_START 129840
<< end >>

